module BCD(
	input[3:0] in_A,
	output reg [6:0] out_B
);

	
always@(*)
begin
	case (in_A)
		4'b0000: out_B = 7'b1000000; // 0 = 0111111
		4'b0001: out_B = 7'b1111001; // 1 = 0000110
		4'b0010: out_B = 7'b0100100; // 2 = 1011011
		4'b0011: out_B = 7'b0110000; // 3 = 1001111
		4'b0100: out_B = 7'b0011001; // 4 = 1100110
		4'b0101: out_B = 7'b0010010; // 5 = 1101101
		4'b0110: out_B = 7'b0000010; // 6 = 1111101
		4'b0111: out_B = 7'b1111000; // 7 = 0000111
		4'b1000: out_B = 7'b0000000; // 8 = 1111111
		4'b1001: out_B = 7'b0010000; // 9 = 1101111
		4'b1010: out_B = 7'b0001000; // A = 1110111
		4'b1011: out_B = 7'b0000011; // B = 1111100
		4'b1100: out_B = 7'b1000110; // C = 0111001
		4'b1101: out_B = 7'b0100001; // D = 1011110
		4'b1110: out_B = 7'b0000110; // E = 1111001
		4'b1111: out_B = 7'b0111111; // - = 1000000
	endcase
end

endmodule
